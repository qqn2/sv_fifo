class generator;

rand transaction trans;

task main();
	trans = new();
	
endtask : main







endclass